module extend(input logic [24:0] imm,
				  input logic [1:0] immsrc,
				  output logic [31:0] immext);
	
	always_comb begin
    case (immsrc)
        2'b00: immext= {{20{imm[24]}},imm[24:13]};												//I type
        2'b01: immext= {{20{imm[24]}},imm[0],imm[23:18],imm[4:1],1'b0}; 				//B type
		  2'b10: immext= {{20{imm[24]}},imm[24:18],imm[4:0]};       				//S type
		  2'b11: immext= {{12{imm[24]}},imm[12:5],imm[13],imm[23:14],1'b0};	//J type
        default: immext = 32'hxxxx_xxxx;
    endcase
	end
	
endmodule
